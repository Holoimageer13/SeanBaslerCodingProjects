CIRCUIT FILE FOR EXP 10-1
VG32 3 2 sin(0,10,200K,0,0,90)
R31 3 1 50
R20 2 0 100
C10 1 0 0.010U IC = 0
.TRAN 0.1E-6 10E-6 0.01E-6 UIC
.PROBE
.END