Name: Sean Basler  Problem:3  Experiment: 3 ;Title
V1 5 0 DC 50 ;Voltage Source
R1 5 4 10	 ; 10 ohm Resistor in circuit
R2 5 2 90	 ; 90 ohm Resistor in circuit
R3 4 6 90	 ; 90 ohm Resistor in dummy node for the dummy voltage 
R4 1 2 30	 ; 30 ohm Resistor in circuit
R5 2 3 30	 ; 30 ohm Resistor in circuit
R6 1 0 10	 ; 10 ohm Resistor in circuit
R7 3 0 90	 ; 90 ohm Resistor in circuit
VD1 6 1 DC 0 ;Dummy used to detect current between 4 and 1
H1 4 3 VD1 30;implementation of current dependent voltage source
.OP
.END